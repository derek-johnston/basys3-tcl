/////////////////////////////////////////////////////////////////////////////////////////
// top.v
// Developed By: 
// Last Modified: 
/////////////////////////////////////////////////////////////////////////////////////////
module top();
endmodule